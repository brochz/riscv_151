
`define RESP_OKAY   0
`define RESP_EXOKAY 1
`define RESP_SLVERR 2
`define RESP_DECERR 3

`define BURST_FIXED 0
`define BURST_INCR  1
`define BURST_WRAP  2

`define LOCK_NORMAL 0
`define LOCK_EXCLSV 1
`define LOCK_LOCKED 2

